
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_fixed_to_float_top.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_fixed_to_float_top.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_fixed_to_float_top.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.grp_convert_ac_fixed_ac_float_25_2_8_0_Pipeline_VITIS_LOOP_213_fu_154.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.grp_convert_ac_fixed_ac_float_25_2_8_0_Pipeline_VITIS_LOOP_213_fu_154.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_fixed_to_float_top.grp_convert_ac_fixed_ac_float_25_2_8_0_s_fu_41.grp_convert_ac_fixed_ac_float_25_2_8_0_Pipeline_VITIS_LOOP_213_fu_154.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;


    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);





    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
